module template (input p62, output p44);
endmodule